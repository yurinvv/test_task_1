package tb_pckg;
	`include "Driver.svh"
	`include "OutData.svh"
	`include "Monitor.svh"
	`include "Scoreboard.svh"
	`include "Environment.svh"
	`include "Test_Check_48.svh"
	`include "Test_Check_1008.svh"
	`include "Test_Check_6144.svh"
endpackage