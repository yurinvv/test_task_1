class OutData;
	bit sov;
	bit [31:0] vector_data;
	bit eov;
endclass